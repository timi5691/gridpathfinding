module update

import mystructs

pub fn update(mut app mystructs.App) {

}